
typedef enum bit {write, read} i2c_op_t;

