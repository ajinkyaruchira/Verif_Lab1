package mypack;

	typedef enum bit {READ = 1'b0 , WRITE = 1'b1} i2c_op_t;
	i2c_op_t op;

endpackage;